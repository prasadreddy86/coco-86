//Fifo design with 16 bit deapth
//***************************************************************************//

module fifo(
             output reg rd_data[n-1:0],
             output reg ful_emptybar,
             output reg             
            );

endmodule
